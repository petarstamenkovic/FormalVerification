
module sv_model(clk, rst, x, y);
  input clk, rst;
  input [1023:0] x;
  output [1023:0] y;
  wire clk, rst;
  wire [1023:0] x;
  wire [1023:0] y;
  wire [7:0] cnt;
  wire n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089;
  wire n_3090, n_3091, n_3093, n_3095, n_3096, n_3098, n_3099, n_3100;
  wire n_3101, n_3102, n_3103, n_3104, n_3105, n_3107, n_3108, n_3109;
  wire n_3110, n_3111, n_3112, n_3114, n_3115, n_3116, n_3118, n_3119;
  wire n_3121, n_3122, n_3124, n_3134, n_3135, n_3138, n_3139, n_3140;
  wire n_3141, n_3142, n_3143, n_3146, n_3149, n_3159, n_3160, n_3161;
  wire n_3164, n_3167, n_3170, n_3173, n_3188, n_3189, n_3190, n_3191;
  wire n_3192, n_3193, n_3194, n_3207, n_3208, n_3209, n_3210, n_3211;
  wire n_3212, n_3215, n_3218, n_3231, n_3232, n_3233, n_3234, n_3235;
  wire n_3236, n_3241, n_3242, n_3245, n_3248, n_3253, n_3254, n_3263;
  wire n_3264, n_3265, n_3266, n_3269, n_3272, n_3277, n_3278, n_3287;
  wire n_3288, n_3289, n_3290, n_3297, n_3298, n_3299, n_3310, n_3311;
  wire n_3312, n_3313, n_3314, n_3331, n_3332, n_3333, n_3334, n_3335;
  wire n_3336, n_3337, n_3338, n_3367, n_3368, n_3369, n_3370, n_3373;
  wire n_3374, n_3375, n_3376, n_3379, n_3381, n_3382, n_3383, n_3384;
  wire n_3385, n_3386;
  assign y[30] = 1'b0;
  assign y[31] = 1'b0;
  assign y[32] = 1'b0;
  assign y[33] = 1'b0;
  assign y[34] = 1'b0;
  assign y[35] = 1'b0;
  assign y[36] = 1'b0;
  assign y[37] = 1'b0;
  assign y[38] = 1'b0;
  assign y[39] = 1'b0;
  assign y[40] = 1'b0;
  assign y[41] = 1'b0;
  assign y[42] = 1'b0;
  assign y[43] = 1'b0;
  assign y[44] = 1'b0;
  assign y[45] = 1'b0;
  assign y[46] = 1'b0;
  assign y[47] = 1'b0;
  assign y[48] = 1'b0;
  assign y[49] = 1'b0;
  assign y[50] = 1'b0;
  assign y[51] = 1'b0;
  assign y[52] = 1'b0;
  assign y[53] = 1'b0;
  assign y[54] = 1'b0;
  assign y[55] = 1'b0;
  assign y[56] = 1'b0;
  assign y[57] = 1'b0;
  assign y[58] = 1'b0;
  assign y[59] = 1'b0;
  assign y[60] = 1'b0;
  assign y[61] = 1'b0;
  assign y[62] = 1'b0;
  assign y[63] = 1'b0;
  assign y[64] = 1'b0;
  assign y[65] = 1'b0;
  assign y[66] = 1'b0;
  assign y[67] = 1'b0;
  assign y[68] = 1'b0;
  assign y[69] = 1'b0;
  assign y[70] = 1'b0;
  assign y[71] = 1'b0;
  assign y[72] = 1'b0;
  assign y[73] = 1'b0;
  assign y[74] = 1'b0;
  assign y[75] = 1'b0;
  assign y[76] = 1'b0;
  assign y[77] = 1'b0;
  assign y[78] = 1'b0;
  assign y[79] = 1'b0;
  assign y[80] = 1'b0;
  assign y[81] = 1'b0;
  assign y[82] = 1'b0;
  assign y[83] = 1'b0;
  assign y[84] = 1'b0;
  assign y[85] = 1'b0;
  assign y[86] = 1'b0;
  assign y[87] = 1'b0;
  assign y[88] = 1'b0;
  assign y[89] = 1'b0;
  assign y[90] = 1'b0;
  assign y[91] = 1'b0;
  assign y[92] = 1'b0;
  assign y[93] = 1'b0;
  assign y[94] = 1'b0;
  assign y[95] = 1'b0;
  assign y[96] = 1'b0;
  assign y[97] = 1'b0;
  assign y[98] = 1'b0;
  assign y[99] = 1'b0;
  assign y[100] = 1'b0;
  assign y[101] = 1'b0;
  assign y[102] = 1'b0;
  assign y[103] = 1'b0;
  assign y[104] = 1'b0;
  assign y[105] = 1'b0;
  assign y[106] = 1'b0;
  assign y[107] = 1'b0;
  assign y[108] = 1'b0;
  assign y[109] = 1'b0;
  assign y[110] = 1'b0;
  assign y[111] = 1'b0;
  assign y[112] = 1'b0;
  assign y[113] = 1'b0;
  assign y[114] = 1'b0;
  assign y[115] = 1'b0;
  assign y[116] = 1'b0;
  assign y[117] = 1'b0;
  assign y[118] = 1'b0;
  assign y[119] = 1'b0;
  assign y[120] = 1'b0;
  assign y[121] = 1'b0;
  assign y[122] = 1'b0;
  assign y[123] = 1'b0;
  assign y[124] = 1'b0;
  assign y[125] = 1'b0;
  assign y[126] = 1'b0;
  assign y[127] = 1'b0;
  assign y[128] = 1'b0;
  assign y[129] = 1'b0;
  assign y[130] = 1'b0;
  assign y[131] = 1'b0;
  assign y[132] = 1'b0;
  assign y[133] = 1'b0;
  assign y[134] = 1'b0;
  assign y[135] = 1'b0;
  assign y[136] = 1'b0;
  assign y[137] = 1'b0;
  assign y[138] = 1'b0;
  assign y[139] = 1'b0;
  assign y[140] = 1'b0;
  assign y[141] = 1'b0;
  assign y[142] = 1'b0;
  assign y[143] = 1'b0;
  assign y[144] = 1'b0;
  assign y[145] = 1'b0;
  assign y[146] = 1'b0;
  assign y[147] = 1'b0;
  assign y[148] = 1'b0;
  assign y[149] = 1'b0;
  assign y[150] = 1'b0;
  assign y[151] = 1'b0;
  assign y[152] = 1'b0;
  assign y[153] = 1'b0;
  assign y[154] = 1'b0;
  assign y[155] = 1'b0;
  assign y[156] = 1'b0;
  assign y[157] = 1'b0;
  assign y[158] = 1'b0;
  assign y[159] = 1'b0;
  assign y[160] = 1'b0;
  assign y[161] = 1'b0;
  assign y[162] = 1'b0;
  assign y[163] = 1'b0;
  assign y[164] = 1'b0;
  assign y[165] = 1'b0;
  assign y[166] = 1'b0;
  assign y[167] = 1'b0;
  assign y[168] = 1'b0;
  assign y[169] = 1'b0;
  assign y[170] = 1'b0;
  assign y[171] = 1'b0;
  assign y[172] = 1'b0;
  assign y[173] = 1'b0;
  assign y[174] = 1'b0;
  assign y[175] = 1'b0;
  assign y[176] = 1'b0;
  assign y[177] = 1'b0;
  assign y[178] = 1'b0;
  assign y[179] = 1'b0;
  assign y[180] = 1'b0;
  assign y[181] = 1'b0;
  assign y[182] = 1'b0;
  assign y[183] = 1'b0;
  assign y[184] = 1'b0;
  assign y[185] = 1'b0;
  assign y[186] = 1'b0;
  assign y[187] = 1'b0;
  assign y[188] = 1'b0;
  assign y[189] = 1'b0;
  assign y[190] = 1'b0;
  assign y[191] = 1'b0;
  assign y[192] = 1'b0;
  assign y[193] = 1'b0;
  assign y[194] = 1'b0;
  assign y[195] = 1'b0;
  assign y[196] = 1'b0;
  assign y[197] = 1'b0;
  assign y[198] = 1'b0;
  assign y[199] = 1'b0;
  assign y[200] = 1'b0;
  assign y[201] = 1'b0;
  assign y[202] = 1'b0;
  assign y[203] = 1'b0;
  assign y[204] = 1'b0;
  assign y[205] = 1'b0;
  assign y[206] = 1'b0;
  assign y[207] = 1'b0;
  assign y[208] = 1'b0;
  assign y[209] = 1'b0;
  assign y[210] = 1'b0;
  assign y[211] = 1'b0;
  assign y[212] = 1'b0;
  assign y[213] = 1'b0;
  assign y[214] = 1'b0;
  assign y[215] = 1'b0;
  assign y[216] = 1'b0;
  assign y[217] = 1'b0;
  assign y[218] = 1'b0;
  assign y[219] = 1'b0;
  assign y[220] = 1'b0;
  assign y[221] = 1'b0;
  assign y[222] = 1'b0;
  assign y[223] = 1'b0;
  assign y[224] = 1'b0;
  assign y[225] = 1'b0;
  assign y[226] = 1'b0;
  assign y[227] = 1'b0;
  assign y[228] = 1'b0;
  assign y[229] = 1'b0;
  assign y[230] = 1'b0;
  assign y[231] = 1'b0;
  assign y[232] = 1'b0;
  assign y[233] = 1'b0;
  assign y[234] = 1'b0;
  assign y[235] = 1'b0;
  assign y[236] = 1'b0;
  assign y[237] = 1'b0;
  assign y[238] = 1'b0;
  assign y[239] = 1'b0;
  assign y[240] = 1'b0;
  assign y[241] = 1'b0;
  assign y[242] = 1'b0;
  assign y[243] = 1'b0;
  assign y[244] = 1'b0;
  assign y[245] = 1'b0;
  assign y[246] = 1'b0;
  assign y[247] = 1'b0;
  assign y[248] = 1'b0;
  assign y[249] = 1'b0;
  assign y[250] = 1'b0;
  assign y[251] = 1'b0;
  assign y[252] = 1'b0;
  assign y[253] = 1'b0;
  assign y[254] = 1'b0;
  assign y[255] = 1'b0;
  assign y[256] = 1'b0;
  assign y[257] = 1'b0;
  assign y[258] = 1'b0;
  assign y[259] = 1'b0;
  assign y[260] = 1'b0;
  assign y[261] = 1'b0;
  assign y[262] = 1'b0;
  assign y[263] = 1'b0;
  assign y[264] = 1'b0;
  assign y[265] = 1'b0;
  assign y[266] = 1'b0;
  assign y[267] = 1'b0;
  assign y[268] = 1'b0;
  assign y[269] = 1'b0;
  assign y[270] = 1'b0;
  assign y[271] = 1'b0;
  assign y[272] = 1'b0;
  assign y[273] = 1'b0;
  assign y[274] = 1'b0;
  assign y[275] = 1'b0;
  assign y[276] = 1'b0;
  assign y[277] = 1'b0;
  assign y[278] = 1'b0;
  assign y[279] = 1'b0;
  assign y[280] = 1'b0;
  assign y[281] = 1'b0;
  assign y[282] = 1'b0;
  assign y[283] = 1'b0;
  assign y[284] = 1'b0;
  assign y[285] = 1'b0;
  assign y[286] = 1'b0;
  assign y[287] = 1'b0;
  assign y[288] = 1'b0;
  assign y[289] = 1'b0;
  assign y[290] = 1'b0;
  assign y[291] = 1'b0;
  assign y[292] = 1'b0;
  assign y[293] = 1'b0;
  assign y[294] = 1'b0;
  assign y[295] = 1'b0;
  assign y[296] = 1'b0;
  assign y[297] = 1'b0;
  assign y[298] = 1'b0;
  assign y[299] = 1'b0;
  assign y[300] = 1'b0;
  assign y[301] = 1'b0;
  assign y[302] = 1'b0;
  assign y[303] = 1'b0;
  assign y[304] = 1'b0;
  assign y[305] = 1'b0;
  assign y[306] = 1'b0;
  assign y[307] = 1'b0;
  assign y[308] = 1'b0;
  assign y[309] = 1'b0;
  assign y[310] = 1'b0;
  assign y[311] = 1'b0;
  assign y[312] = 1'b0;
  assign y[313] = 1'b0;
  assign y[314] = 1'b0;
  assign y[315] = 1'b0;
  assign y[316] = 1'b0;
  assign y[317] = 1'b0;
  assign y[318] = 1'b0;
  assign y[319] = 1'b0;
  assign y[320] = 1'b0;
  assign y[321] = 1'b0;
  assign y[322] = 1'b0;
  assign y[323] = 1'b0;
  assign y[324] = 1'b0;
  assign y[325] = 1'b0;
  assign y[326] = 1'b0;
  assign y[327] = 1'b0;
  assign y[328] = 1'b0;
  assign y[329] = 1'b0;
  assign y[330] = 1'b0;
  assign y[331] = 1'b0;
  assign y[332] = 1'b0;
  assign y[333] = 1'b0;
  assign y[334] = 1'b0;
  assign y[335] = 1'b0;
  assign y[336] = 1'b0;
  assign y[337] = 1'b0;
  assign y[338] = 1'b0;
  assign y[339] = 1'b0;
  assign y[340] = 1'b0;
  assign y[341] = 1'b0;
  assign y[342] = 1'b0;
  assign y[343] = 1'b0;
  assign y[344] = 1'b0;
  assign y[345] = 1'b0;
  assign y[346] = 1'b0;
  assign y[347] = 1'b0;
  assign y[348] = 1'b0;
  assign y[349] = 1'b0;
  assign y[350] = 1'b0;
  assign y[351] = 1'b0;
  assign y[352] = 1'b0;
  assign y[353] = 1'b0;
  assign y[354] = 1'b0;
  assign y[355] = 1'b0;
  assign y[356] = 1'b0;
  assign y[357] = 1'b0;
  assign y[358] = 1'b0;
  assign y[359] = 1'b0;
  assign y[360] = 1'b0;
  assign y[361] = 1'b0;
  assign y[362] = 1'b0;
  assign y[363] = 1'b0;
  assign y[364] = 1'b0;
  assign y[365] = 1'b0;
  assign y[366] = 1'b0;
  assign y[367] = 1'b0;
  assign y[368] = 1'b0;
  assign y[369] = 1'b0;
  assign y[370] = 1'b0;
  assign y[371] = 1'b0;
  assign y[372] = 1'b0;
  assign y[373] = 1'b0;
  assign y[374] = 1'b0;
  assign y[375] = 1'b0;
  assign y[376] = 1'b0;
  assign y[377] = 1'b0;
  assign y[378] = 1'b0;
  assign y[379] = 1'b0;
  assign y[380] = 1'b0;
  assign y[381] = 1'b0;
  assign y[382] = 1'b0;
  assign y[383] = 1'b0;
  assign y[384] = 1'b0;
  assign y[385] = 1'b0;
  assign y[386] = 1'b0;
  assign y[387] = 1'b0;
  assign y[388] = 1'b0;
  assign y[389] = 1'b0;
  assign y[390] = 1'b0;
  assign y[391] = 1'b0;
  assign y[392] = 1'b0;
  assign y[393] = 1'b0;
  assign y[394] = 1'b0;
  assign y[395] = 1'b0;
  assign y[396] = 1'b0;
  assign y[397] = 1'b0;
  assign y[398] = 1'b0;
  assign y[399] = 1'b0;
  assign y[400] = 1'b0;
  assign y[401] = 1'b0;
  assign y[402] = 1'b0;
  assign y[403] = 1'b0;
  assign y[404] = 1'b0;
  assign y[405] = 1'b0;
  assign y[406] = 1'b0;
  assign y[407] = 1'b0;
  assign y[408] = 1'b0;
  assign y[409] = 1'b0;
  assign y[410] = 1'b0;
  assign y[411] = 1'b0;
  assign y[412] = 1'b0;
  assign y[413] = 1'b0;
  assign y[414] = 1'b0;
  assign y[415] = 1'b0;
  assign y[416] = 1'b0;
  assign y[417] = 1'b0;
  assign y[418] = 1'b0;
  assign y[419] = 1'b0;
  assign y[420] = 1'b0;
  assign y[421] = 1'b0;
  assign y[422] = 1'b0;
  assign y[423] = 1'b0;
  assign y[424] = 1'b0;
  assign y[425] = 1'b0;
  assign y[426] = 1'b0;
  assign y[427] = 1'b0;
  assign y[428] = 1'b0;
  assign y[429] = 1'b0;
  assign y[430] = 1'b0;
  assign y[431] = 1'b0;
  assign y[432] = 1'b0;
  assign y[433] = 1'b0;
  assign y[434] = 1'b0;
  assign y[435] = 1'b0;
  assign y[436] = 1'b0;
  assign y[437] = 1'b0;
  assign y[438] = 1'b0;
  assign y[439] = 1'b0;
  assign y[440] = 1'b0;
  assign y[441] = 1'b0;
  assign y[442] = 1'b0;
  assign y[443] = 1'b0;
  assign y[444] = 1'b0;
  assign y[445] = 1'b0;
  assign y[446] = 1'b0;
  assign y[447] = 1'b0;
  assign y[448] = 1'b0;
  assign y[449] = 1'b0;
  assign y[450] = 1'b0;
  assign y[451] = 1'b0;
  assign y[452] = 1'b0;
  assign y[453] = 1'b0;
  assign y[454] = 1'b0;
  assign y[455] = 1'b0;
  assign y[456] = 1'b0;
  assign y[457] = 1'b0;
  assign y[458] = 1'b0;
  assign y[459] = 1'b0;
  assign y[460] = 1'b0;
  assign y[461] = 1'b0;
  assign y[462] = 1'b0;
  assign y[463] = 1'b0;
  assign y[464] = 1'b0;
  assign y[465] = 1'b0;
  assign y[466] = 1'b0;
  assign y[467] = 1'b0;
  assign y[468] = 1'b0;
  assign y[469] = 1'b0;
  assign y[470] = 1'b0;
  assign y[471] = 1'b0;
  assign y[472] = 1'b0;
  assign y[473] = 1'b0;
  assign y[474] = 1'b0;
  assign y[475] = 1'b0;
  assign y[476] = 1'b0;
  assign y[477] = 1'b0;
  assign y[478] = 1'b0;
  assign y[479] = 1'b0;
  assign y[480] = 1'b0;
  assign y[481] = 1'b0;
  assign y[482] = 1'b0;
  assign y[483] = 1'b0;
  assign y[484] = 1'b0;
  assign y[485] = 1'b0;
  assign y[486] = 1'b0;
  assign y[487] = 1'b0;
  assign y[488] = 1'b0;
  assign y[489] = 1'b0;
  assign y[490] = 1'b0;
  assign y[491] = 1'b0;
  assign y[492] = 1'b0;
  assign y[493] = 1'b0;
  assign y[494] = 1'b0;
  assign y[495] = 1'b0;
  assign y[496] = 1'b0;
  assign y[497] = 1'b0;
  assign y[498] = 1'b0;
  assign y[499] = 1'b0;
  assign y[500] = 1'b0;
  assign y[501] = 1'b0;
  assign y[502] = 1'b0;
  assign y[503] = 1'b0;
  assign y[504] = 1'b0;
  assign y[505] = 1'b0;
  assign y[506] = 1'b0;
  assign y[507] = 1'b0;
  assign y[508] = 1'b0;
  assign y[509] = 1'b0;
  assign y[510] = 1'b0;
  assign y[511] = 1'b0;
  assign y[512] = 1'b0;
  assign y[513] = 1'b0;
  assign y[514] = 1'b0;
  assign y[515] = 1'b0;
  assign y[516] = 1'b0;
  assign y[517] = 1'b0;
  assign y[518] = 1'b0;
  assign y[519] = 1'b0;
  assign y[520] = 1'b0;
  assign y[521] = 1'b0;
  assign y[522] = 1'b0;
  assign y[523] = 1'b0;
  assign y[524] = 1'b0;
  assign y[525] = 1'b0;
  assign y[526] = 1'b0;
  assign y[527] = 1'b0;
  assign y[528] = 1'b0;
  assign y[529] = 1'b0;
  assign y[530] = 1'b0;
  assign y[531] = 1'b0;
  assign y[532] = 1'b0;
  assign y[533] = 1'b0;
  assign y[534] = 1'b0;
  assign y[535] = 1'b0;
  assign y[536] = 1'b0;
  assign y[537] = 1'b0;
  assign y[538] = 1'b0;
  assign y[539] = 1'b0;
  assign y[540] = 1'b0;
  assign y[541] = 1'b0;
  assign y[542] = 1'b0;
  assign y[543] = 1'b0;
  assign y[544] = 1'b0;
  assign y[545] = 1'b0;
  assign y[546] = 1'b0;
  assign y[547] = 1'b0;
  assign y[548] = 1'b0;
  assign y[549] = 1'b0;
  assign y[550] = 1'b0;
  assign y[551] = 1'b0;
  assign y[552] = 1'b0;
  assign y[553] = 1'b0;
  assign y[554] = 1'b0;
  assign y[555] = 1'b0;
  assign y[556] = 1'b0;
  assign y[557] = 1'b0;
  assign y[558] = 1'b0;
  assign y[559] = 1'b0;
  assign y[560] = 1'b0;
  assign y[561] = 1'b0;
  assign y[562] = 1'b0;
  assign y[563] = 1'b0;
  assign y[564] = 1'b0;
  assign y[565] = 1'b0;
  assign y[566] = 1'b0;
  assign y[567] = 1'b0;
  assign y[568] = 1'b0;
  assign y[569] = 1'b0;
  assign y[570] = 1'b0;
  assign y[571] = 1'b0;
  assign y[572] = 1'b0;
  assign y[573] = 1'b0;
  assign y[574] = 1'b0;
  assign y[575] = 1'b0;
  assign y[576] = 1'b0;
  assign y[577] = 1'b0;
  assign y[578] = 1'b0;
  assign y[579] = 1'b0;
  assign y[580] = 1'b0;
  assign y[581] = 1'b0;
  assign y[582] = 1'b0;
  assign y[583] = 1'b0;
  assign y[584] = 1'b0;
  assign y[585] = 1'b0;
  assign y[586] = 1'b0;
  assign y[587] = 1'b0;
  assign y[588] = 1'b0;
  assign y[589] = 1'b0;
  assign y[590] = 1'b0;
  assign y[591] = 1'b0;
  assign y[592] = 1'b0;
  assign y[593] = 1'b0;
  assign y[594] = 1'b0;
  assign y[595] = 1'b0;
  assign y[596] = 1'b0;
  assign y[597] = 1'b0;
  assign y[598] = 1'b0;
  assign y[599] = 1'b0;
  assign y[600] = 1'b0;
  assign y[601] = 1'b0;
  assign y[602] = 1'b0;
  assign y[603] = 1'b0;
  assign y[604] = 1'b0;
  assign y[605] = 1'b0;
  assign y[606] = 1'b0;
  assign y[607] = 1'b0;
  assign y[608] = 1'b0;
  assign y[609] = 1'b0;
  assign y[610] = 1'b0;
  assign y[611] = 1'b0;
  assign y[612] = 1'b0;
  assign y[613] = 1'b0;
  assign y[614] = 1'b0;
  assign y[615] = 1'b0;
  assign y[616] = 1'b0;
  assign y[617] = 1'b0;
  assign y[618] = 1'b0;
  assign y[619] = 1'b0;
  assign y[620] = 1'b0;
  assign y[621] = 1'b0;
  assign y[622] = 1'b0;
  assign y[623] = 1'b0;
  assign y[624] = 1'b0;
  assign y[625] = 1'b0;
  assign y[626] = 1'b0;
  assign y[627] = 1'b0;
  assign y[628] = 1'b0;
  assign y[629] = 1'b0;
  assign y[630] = 1'b0;
  assign y[631] = 1'b0;
  assign y[632] = 1'b0;
  assign y[633] = 1'b0;
  assign y[634] = 1'b0;
  assign y[635] = 1'b0;
  assign y[636] = 1'b0;
  assign y[637] = 1'b0;
  assign y[638] = 1'b0;
  assign y[639] = 1'b0;
  assign y[640] = 1'b0;
  assign y[641] = 1'b0;
  assign y[642] = 1'b0;
  assign y[643] = 1'b0;
  assign y[644] = 1'b0;
  assign y[645] = 1'b0;
  assign y[646] = 1'b0;
  assign y[647] = 1'b0;
  assign y[648] = 1'b0;
  assign y[649] = 1'b0;
  assign y[650] = 1'b0;
  assign y[651] = 1'b0;
  assign y[652] = 1'b0;
  assign y[653] = 1'b0;
  assign y[654] = 1'b0;
  assign y[655] = 1'b0;
  assign y[656] = 1'b0;
  assign y[657] = 1'b0;
  assign y[658] = 1'b0;
  assign y[659] = 1'b0;
  assign y[660] = 1'b0;
  assign y[661] = 1'b0;
  assign y[662] = 1'b0;
  assign y[663] = 1'b0;
  assign y[664] = 1'b0;
  assign y[665] = 1'b0;
  assign y[666] = 1'b0;
  assign y[667] = 1'b0;
  assign y[668] = 1'b0;
  assign y[669] = 1'b0;
  assign y[670] = 1'b0;
  assign y[671] = 1'b0;
  assign y[672] = 1'b0;
  assign y[673] = 1'b0;
  assign y[674] = 1'b0;
  assign y[675] = 1'b0;
  assign y[676] = 1'b0;
  assign y[677] = 1'b0;
  assign y[678] = 1'b0;
  assign y[679] = 1'b0;
  assign y[680] = 1'b0;
  assign y[681] = 1'b0;
  assign y[682] = 1'b0;
  assign y[683] = 1'b0;
  assign y[684] = 1'b0;
  assign y[685] = 1'b0;
  assign y[686] = 1'b0;
  assign y[687] = 1'b0;
  assign y[688] = 1'b0;
  assign y[689] = 1'b0;
  assign y[690] = 1'b0;
  assign y[691] = 1'b0;
  assign y[692] = 1'b0;
  assign y[693] = 1'b0;
  assign y[694] = 1'b0;
  assign y[695] = 1'b0;
  assign y[696] = 1'b0;
  assign y[697] = 1'b0;
  assign y[698] = 1'b0;
  assign y[699] = 1'b0;
  assign y[700] = 1'b0;
  assign y[701] = 1'b0;
  assign y[702] = 1'b0;
  assign y[703] = 1'b0;
  assign y[704] = 1'b0;
  assign y[705] = 1'b0;
  assign y[706] = 1'b0;
  assign y[707] = 1'b0;
  assign y[708] = 1'b0;
  assign y[709] = 1'b0;
  assign y[710] = 1'b0;
  assign y[711] = 1'b0;
  assign y[712] = 1'b0;
  assign y[713] = 1'b0;
  assign y[714] = 1'b0;
  assign y[715] = 1'b0;
  assign y[716] = 1'b0;
  assign y[717] = 1'b0;
  assign y[718] = 1'b0;
  assign y[719] = 1'b0;
  assign y[720] = 1'b0;
  assign y[721] = 1'b0;
  assign y[722] = 1'b0;
  assign y[723] = 1'b0;
  assign y[724] = 1'b0;
  assign y[725] = 1'b0;
  assign y[726] = 1'b0;
  assign y[727] = 1'b0;
  assign y[728] = 1'b0;
  assign y[729] = 1'b0;
  assign y[730] = 1'b0;
  assign y[731] = 1'b0;
  assign y[732] = 1'b0;
  assign y[733] = 1'b0;
  assign y[734] = 1'b0;
  assign y[735] = 1'b0;
  assign y[736] = 1'b0;
  assign y[737] = 1'b0;
  assign y[738] = 1'b0;
  assign y[739] = 1'b0;
  assign y[740] = 1'b0;
  assign y[741] = 1'b0;
  assign y[742] = 1'b0;
  assign y[743] = 1'b0;
  assign y[744] = 1'b0;
  assign y[745] = 1'b0;
  assign y[746] = 1'b0;
  assign y[747] = 1'b0;
  assign y[748] = 1'b0;
  assign y[749] = 1'b0;
  assign y[750] = 1'b0;
  assign y[751] = 1'b0;
  assign y[752] = 1'b0;
  assign y[753] = 1'b0;
  assign y[754] = 1'b0;
  assign y[755] = 1'b0;
  assign y[756] = 1'b0;
  assign y[757] = 1'b0;
  assign y[758] = 1'b0;
  assign y[759] = 1'b0;
  assign y[760] = 1'b0;
  assign y[761] = 1'b0;
  assign y[762] = 1'b0;
  assign y[763] = 1'b0;
  assign y[764] = 1'b0;
  assign y[765] = 1'b0;
  assign y[766] = 1'b0;
  assign y[767] = 1'b0;
  assign y[768] = 1'b0;
  assign y[769] = 1'b0;
  assign y[770] = 1'b0;
  assign y[771] = 1'b0;
  assign y[772] = 1'b0;
  assign y[773] = 1'b0;
  assign y[774] = 1'b0;
  assign y[775] = 1'b0;
  assign y[776] = 1'b0;
  assign y[777] = 1'b0;
  assign y[778] = 1'b0;
  assign y[779] = 1'b0;
  assign y[780] = 1'b0;
  assign y[781] = 1'b0;
  assign y[782] = 1'b0;
  assign y[783] = 1'b0;
  assign y[784] = 1'b0;
  assign y[785] = 1'b0;
  assign y[786] = 1'b0;
  assign y[787] = 1'b0;
  assign y[788] = 1'b0;
  assign y[789] = 1'b0;
  assign y[790] = 1'b0;
  assign y[791] = 1'b0;
  assign y[792] = 1'b0;
  assign y[793] = 1'b0;
  assign y[794] = 1'b0;
  assign y[795] = 1'b0;
  assign y[796] = 1'b0;
  assign y[797] = 1'b0;
  assign y[798] = 1'b0;
  assign y[799] = 1'b0;
  assign y[800] = 1'b0;
  assign y[801] = 1'b0;
  assign y[802] = 1'b0;
  assign y[803] = 1'b0;
  assign y[804] = 1'b0;
  assign y[805] = 1'b0;
  assign y[806] = 1'b0;
  assign y[807] = 1'b0;
  assign y[808] = 1'b0;
  assign y[809] = 1'b0;
  assign y[810] = 1'b0;
  assign y[811] = 1'b0;
  assign y[812] = 1'b0;
  assign y[813] = 1'b0;
  assign y[814] = 1'b0;
  assign y[815] = 1'b0;
  assign y[816] = 1'b0;
  assign y[817] = 1'b0;
  assign y[818] = 1'b0;
  assign y[819] = 1'b0;
  assign y[820] = 1'b0;
  assign y[821] = 1'b0;
  assign y[822] = 1'b0;
  assign y[823] = 1'b0;
  assign y[824] = 1'b0;
  assign y[825] = 1'b0;
  assign y[826] = 1'b0;
  assign y[827] = 1'b0;
  assign y[828] = 1'b0;
  assign y[829] = 1'b0;
  assign y[830] = 1'b0;
  assign y[831] = 1'b0;
  assign y[832] = 1'b0;
  assign y[833] = 1'b0;
  assign y[834] = 1'b0;
  assign y[835] = 1'b0;
  assign y[836] = 1'b0;
  assign y[837] = 1'b0;
  assign y[838] = 1'b0;
  assign y[839] = 1'b0;
  assign y[840] = 1'b0;
  assign y[841] = 1'b0;
  assign y[842] = 1'b0;
  assign y[843] = 1'b0;
  assign y[844] = 1'b0;
  assign y[845] = 1'b0;
  assign y[846] = 1'b0;
  assign y[847] = 1'b0;
  assign y[848] = 1'b0;
  assign y[849] = 1'b0;
  assign y[850] = 1'b0;
  assign y[851] = 1'b0;
  assign y[852] = 1'b0;
  assign y[853] = 1'b0;
  assign y[854] = 1'b0;
  assign y[855] = 1'b0;
  assign y[856] = 1'b0;
  assign y[857] = 1'b0;
  assign y[858] = 1'b0;
  assign y[859] = 1'b0;
  assign y[860] = 1'b0;
  assign y[861] = 1'b0;
  assign y[862] = 1'b0;
  assign y[863] = 1'b0;
  assign y[864] = 1'b0;
  assign y[865] = 1'b0;
  assign y[866] = 1'b0;
  assign y[867] = 1'b0;
  assign y[868] = 1'b0;
  assign y[869] = 1'b0;
  assign y[870] = 1'b0;
  assign y[871] = 1'b0;
  assign y[872] = 1'b0;
  assign y[873] = 1'b0;
  assign y[874] = 1'b0;
  assign y[875] = 1'b0;
  assign y[876] = 1'b0;
  assign y[877] = 1'b0;
  assign y[878] = 1'b0;
  assign y[879] = 1'b0;
  assign y[880] = 1'b0;
  assign y[881] = 1'b0;
  assign y[882] = 1'b0;
  assign y[883] = 1'b0;
  assign y[884] = 1'b0;
  assign y[885] = 1'b0;
  assign y[886] = 1'b0;
  assign y[887] = 1'b0;
  assign y[888] = 1'b0;
  assign y[889] = 1'b0;
  assign y[890] = 1'b0;
  assign y[891] = 1'b0;
  assign y[892] = 1'b0;
  assign y[893] = 1'b0;
  assign y[894] = 1'b0;
  assign y[895] = 1'b0;
  assign y[896] = 1'b0;
  assign y[897] = 1'b0;
  assign y[898] = 1'b0;
  assign y[899] = 1'b0;
  assign y[900] = 1'b0;
  assign y[901] = 1'b0;
  assign y[902] = 1'b0;
  assign y[903] = 1'b0;
  assign y[904] = 1'b0;
  assign y[905] = 1'b0;
  assign y[906] = 1'b0;
  assign y[907] = 1'b0;
  assign y[908] = 1'b0;
  assign y[909] = 1'b0;
  assign y[910] = 1'b0;
  assign y[911] = 1'b0;
  assign y[912] = 1'b0;
  assign y[913] = 1'b0;
  assign y[914] = 1'b0;
  assign y[915] = 1'b0;
  assign y[916] = 1'b0;
  assign y[917] = 1'b0;
  assign y[918] = 1'b0;
  assign y[919] = 1'b0;
  assign y[920] = 1'b0;
  assign y[921] = 1'b0;
  assign y[922] = 1'b0;
  assign y[923] = 1'b0;
  assign y[924] = 1'b0;
  assign y[925] = 1'b0;
  assign y[926] = 1'b0;
  assign y[927] = 1'b0;
  assign y[928] = 1'b0;
  assign y[929] = 1'b0;
  assign y[930] = 1'b0;
  assign y[931] = 1'b0;
  assign y[932] = 1'b0;
  assign y[933] = 1'b0;
  assign y[934] = 1'b0;
  assign y[935] = 1'b0;
  assign y[936] = 1'b0;
  assign y[937] = 1'b0;
  assign y[938] = 1'b0;
  assign y[939] = 1'b0;
  assign y[940] = 1'b0;
  assign y[941] = 1'b0;
  assign y[942] = 1'b0;
  assign y[943] = 1'b0;
  assign y[944] = 1'b0;
  assign y[945] = 1'b0;
  assign y[946] = 1'b0;
  assign y[947] = 1'b0;
  assign y[948] = 1'b0;
  assign y[949] = 1'b0;
  assign y[950] = 1'b0;
  assign y[951] = 1'b0;
  assign y[952] = 1'b0;
  assign y[953] = 1'b0;
  assign y[954] = 1'b0;
  assign y[955] = 1'b0;
  assign y[956] = 1'b0;
  assign y[957] = 1'b0;
  assign y[958] = 1'b0;
  assign y[959] = 1'b0;
  assign y[960] = 1'b0;
  assign y[961] = 1'b0;
  assign y[962] = 1'b0;
  assign y[963] = 1'b0;
  assign y[964] = 1'b0;
  assign y[965] = 1'b0;
  assign y[966] = 1'b0;
  assign y[967] = 1'b0;
  assign y[968] = 1'b0;
  assign y[969] = 1'b0;
  assign y[970] = 1'b0;
  assign y[971] = 1'b0;
  assign y[972] = 1'b0;
  assign y[973] = 1'b0;
  assign y[974] = 1'b0;
  assign y[975] = 1'b0;
  assign y[976] = 1'b0;
  assign y[977] = 1'b0;
  assign y[978] = 1'b0;
  assign y[979] = 1'b0;
  assign y[980] = 1'b0;
  assign y[981] = 1'b0;
  assign y[982] = 1'b0;
  assign y[983] = 1'b0;
  assign y[984] = 1'b0;
  assign y[985] = 1'b0;
  assign y[986] = 1'b0;
  assign y[987] = 1'b0;
  assign y[988] = 1'b0;
  assign y[989] = 1'b0;
  assign y[990] = 1'b0;
  assign y[991] = 1'b0;
  assign y[992] = 1'b0;
  assign y[993] = 1'b0;
  assign y[994] = 1'b0;
  assign y[995] = 1'b0;
  assign y[996] = 1'b0;
  assign y[997] = 1'b0;
  assign y[998] = 1'b0;
  assign y[999] = 1'b0;
  assign y[1000] = 1'b0;
  assign y[1001] = 1'b0;
  assign y[1002] = 1'b0;
  assign y[1003] = 1'b0;
  assign y[1004] = 1'b0;
  assign y[1005] = 1'b0;
  assign y[1006] = 1'b0;
  assign y[1007] = 1'b0;
  assign y[1008] = 1'b0;
  assign y[1009] = 1'b0;
  assign y[1010] = 1'b0;
  assign y[1011] = 1'b0;
  assign y[1012] = 1'b0;
  assign y[1013] = 1'b0;
  assign y[1014] = 1'b0;
  assign y[1015] = 1'b0;
  assign y[1016] = 1'b0;
  assign y[1017] = 1'b0;
  assign y[1018] = 1'b0;
  assign y[1019] = 1'b0;
  assign y[1020] = 1'b0;
  assign y[1021] = 1'b0;
  assign y[1022] = 1'b0;
  assign y[1023] = 1'b0;
  CDN_flop \cnt_reg[0] (.clk (clk), .d (n_3085), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[0]));
  CDN_flop \cnt_reg[1] (.clk (clk), .d (n_3112), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[1]));
  CDN_flop \cnt_reg[2] (.clk (clk), .d (n_3098), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[2]));
  CDN_flop \cnt_reg[3] (.clk (clk), .d (n_3107), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[3]));
  CDN_flop \cnt_reg[4] (.clk (clk), .d (n_3100), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[4]));
  CDN_flop \cnt_reg[5] (.clk (clk), .d (n_3108), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[5]));
  CDN_flop \cnt_reg[6] (.clk (clk), .d (n_3103), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[6]));
  CDN_flop \cnt_reg[7] (.clk (clk), .d (n_3110), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (cnt[7]));
  or g15 (n_3099, n_3095, n_3096);
  or g43 (n_3088, cnt[6], cnt[7]);
  or g44 (n_3089, cnt[5], n_3088);
  or g46 (n_3122, n_3089, n_3121);
  nand g1020 (n_3096, cnt[2], cnt[3]);
  or g1023 (n_3121, wc, cnt[3]);
  not gc (wc, cnt[4]);
  or g1025 (n_3105, n_3088, wc0);
  not gc0 (wc0, cnt[5]);
  or g1226 (n_3109, wc1, n_3102);
  not gc1 (wc1, cnt[6]);
  or g1259 (n_3101, n_3099, wc2);
  not gc2 (wc2, cnt[4]);
  or g1262 (n_3102, n_3101, wc3);
  not gc3 (wc3, cnt[5]);
  not g1457 (n_3085, cnt[0]);
  not g1458 (n_3086, rst);
  or g1462 (n_3093, cnt[0], cnt[1]);
  nand g1463 (n_3095, cnt[0], cnt[1]);
  or g1503 (n_3142, cnt[1], wc4);
  not gc4 (wc4, cnt[2]);
  or g1662 (y[0], wc5, n_3314);
  not gc5 (wc5, n_3242);
  or g1663 (y[1], n_3266, wc6);
  not gc6 (wc6, y[11]);
  or g1664 (n_3314, wc7, n_3313);
  not gc7 (wc7, n_3312);
  or g1665 (y[13], n_3337, n_3338);
  or g1666 (y[14], n_3088, n_3194);
  nand g1667 (n_3266, n_3264, n_3265);
  or g1668 (y[3], n_3236, wc8);
  not gc8 (wc8, n_3235);
  or g1669 (n_3118, rst, wc9);
  not gc9 (wc9, n_3272);
  nand g1670 (y[16], n_3277, n_3278);
  or g1671 (y[8], wc10, n_3299);
  not gc10 (wc10, n_3119);
  nand g1672 (y[12], n_3289, n_3290);
  nand g1673 (n_3313, n_3310, n_3311);
  nand g1674 (n_3337, n_3333, n_3334);
  or g1675 (y[9], n_3212, wc11);
  not gc11 (wc11, n_3096);
  or g1676 (n_3194, n_3192, n_3193);
  nand g1677 (n_3334, cnt[1], n_3135);
  or g1678 (n_3289, cnt[1], wc12);
  not gc12 (wc12, n_3135);
  nand g1679 (n_3338, n_3335, n_3336);
  or g1680 (n_3265, cnt[2], n_3263);
  or g1681 (n_3277, wc13, n_3119);
  not gc13 (wc13, cnt[2]);
  or g1682 (n_3311, cnt[2], n_3119);
  nand g1685 (n_3299, n_3297, n_3298);
  or g1686 (n_3272, wc14, n_3109);
  not gc14 (wc14, cnt[7]);
  nand g1687 (n_3367, n_3109, cnt[7]);
  or g1688 (n_3368, n_3109, cnt[7]);
  nand g1689 (n_3110, n_3367, n_3368);
  nand g1690 (y[10], n_3253, n_3254);
  nand g1691 (n_3236, n_3233, n_3234);
  or g1692 (n_3212, n_3089, n_3211);
  or g1693 (n_3119, cnt[3], n_3091);
  nand g1694 (n_3192, n_3188, n_3189);
  or g1695 (n_3211, wc15, n_3210);
  not gc15 (wc15, n_3209);
  or g1696 (n_3335, n_3331, wc16);
  not gc16 (wc16, cnt[2]);
  or g1697 (n_3235, cnt[2], n_3232);
  nand g1698 (n_3369, cnt[6], n_3102);
  or g1699 (n_3370, cnt[6], n_3102);
  nand g1700 (n_3103, n_3369, n_3370);
  or g1701 (n_3310, n_3111, n_3114);
  or g1702 (n_3234, cnt[3], n_3231);
  or g1703 (n_3297, wc17, n_3115);
  not gc17 (wc17, n_3139);
  or g1704 (n_3336, n_3093, n_3332);
  or g1705 (n_3290, cnt[2], n_3288);
  nand g1706 (y[15], n_3241, n_3242);
  or g1709 (n_3278, n_3091, n_3104);
  or g1710 (n_3245, y[29], wc18);
  not gc18 (wc18, n_3138);
  nand g1711 (n_3135, n_3269, n_3114);
  or g1712 (n_3253, n_3115, n_3116);
  or g1713 (n_3107, wc19, n_3161);
  not gc19 (wc19, n_3104);
  or g1714 (y[11], cnt[2], n_3248);
  or g1717 (n_3263, n_3115, n_3111);
  or g1718 (n_3264, n_3095, n_3114);
  or g1719 (n_3254, cnt[1], n_3114);
  or g1720 (n_3248, n_3122, n_3093);
  or g1721 (n_3269, wc20, n_3122);
  not gc20 (wc20, cnt[2]);
  or g1722 (n_3138, cnt[4], n_3173);
  or g1723 (n_3232, wc21, n_3122);
  not gc21 (wc21, n_3093);
  or g1724 (n_3242, n_3090, n_3099);
  or g1725 (n_3241, n_3105, n_3134);
  or g1726 (n_3288, n_3287, wc22);
  not gc22 (wc22, cnt[1]);
  or g1727 (n_3231, n_3089, wc23);
  not gc23 (wc23, n_3124);
  or g1728 (n_3233, n_3090, n_3116);
  or g1729 (n_3218, wc24, n_3090);
  not gc24 (wc24, n_3096);
  or g1730 (n_3298, n_3122, wc25);
  not gc25 (wc25, n_3124);
  or g1731 (n_3312, n_3116, n_3122);
  nand g1732 (n_3373, n_3101, cnt[5]);
  or g1733 (n_3374, n_3101, cnt[5]);
  nand g1734 (n_3108, n_3373, n_3374);
  or g1735 (n_3332, n_3090, n_3096);
  nand g1736 (n_3210, n_3207, n_3208);
  or g1737 (n_3333, n_3089, n_3134);
  or g1738 (n_3114, n_3090, n_3104);
  or g1739 (n_3115, cnt[3], n_3090);
  nand g1740 (n_3193, n_3190, n_3191);
  or g1741 (n_3331, n_3287, wc26);
  not gc26 (wc26, n_3095);
  or g1742 (n_3091, n_3087, n_3090);
  nand g1743 (n_3161, n_3159, n_3160);
  or g1744 (n_3188, cnt[4], wc27);
  not gc27 (wc27, n_3140);
  or g1745 (n_3134, n_3170, wc28);
  not gc28 (wc28, cnt[4]);
  nand g1746 (n_3124, n_3116, n_3215);
  or g1747 (n_3140, cnt[5], wc29);
  not gc29 (wc29, n_3167);
  or g1748 (n_3287, n_3121, n_3105);
  nand g1749 (n_3375, cnt[4], n_3099);
  or g1750 (n_3376, cnt[4], n_3099);
  nand g1751 (n_3100, n_3375, n_3376);
  or g1752 (n_3159, cnt[3], n_3190);
  or g1753 (n_3207, cnt[3], wc30);
  not gc30 (wc30, n_3143);
  or g1754 (n_3090, cnt[4], n_3089);
  nand g1755 (n_3191, n_3141, cnt[4]);
  or g1756 (n_3173, n_3105, n_3096);
  or g1757 (n_3170, n_3093, n_3104);
  nand g1758 (n_3167, cnt[2], n_3093);
  nand g1759 (n_3139, n_3111, n_3164);
  nand g1760 (n_3112, n_3087, n_3111);
  nand g1761 (n_3209, cnt[3], n_3093);
  or g1762 (n_3190, wc31, n_3095);
  not gc31 (wc31, cnt[2]);
  nand g1763 (n_3160, cnt[3], n_3095);
  nand g1764 (n_3143, cnt[0], n_3149);
  or g1765 (n_3141, cnt[3], wc32);
  not gc32 (wc32, n_3146);
  or g1768 (n_3215, cnt[2], n_3095);
  or g1769 (n_3116, wc33, n_3093);
  not gc33 (wc33, cnt[2]);
  nand g1770 (n_3208, n_3142, cnt[4]);
  nand g1773 (n_3379, cnt[2], n_3095);
  nand g1775 (n_3098, n_3379, n_3215);
  nand g1776 (n_3164, cnt[1], cnt[2]);
  or g1777 (n_3381, wc34, y[25]);
  not gc34 (wc34, y[17]);
  or g1778 (n_3382, y[17], wc35);
  not gc35 (wc35, y[25]);
  nand g1779 (n_3083, n_3381, n_3382);
  or g1780 (n_3149, cnt[4], cnt[1]);
  or g1781 (n_3146, cnt[1], cnt[2]);
  or g1782 (n_3189, cnt[3], cnt[5]);
  or g1783 (n_3383, wc36, y[28]);
  not gc36 (wc36, y[17]);
  or g1784 (n_3384, y[17], wc37);
  not gc37 (wc37, y[28]);
  nand g1785 (n_3084, n_3383, n_3384);
  or g1786 (n_3104, cnt[2], wc38);
  not gc38 (wc38, cnt[3]);
  or g1787 (n_3385, wc39, y[23]);
  not gc39 (wc39, y[17]);
  or g1788 (n_3386, y[17], wc40);
  not gc40 (wc40, y[23]);
  nand g1789 (n_3082, n_3385, n_3386);
  or g1790 (n_3087, wc41, cnt[1]);
  not gc41 (wc41, cnt[0]);
  or g1791 (n_3111, cnt[0], wc42);
  not gc42 (wc42, cnt[1]);
  nor g1792 (y[2], y[29], n_3093);
  nor g1793 (y[5], y[29], n_3087);
  and g1794 (y[4], wc43, cnt[2]);
  not gc43 (wc43, n_3091);
  nor g1795 (y[7], n_3095, n_3218);
  nor g1796 (y[6], n_3245, n_3111);
  CDN_flop \lfsr_reg[0] (.clk (clk), .d (y[18]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b1), .q (y[17]));
  CDN_flop \lfsr_reg[1] (.clk (clk), .d (y[19]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[18]));
  CDN_flop \lfsr_reg[2] (.clk (clk), .d (y[20]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[19]));
  CDN_flop \lfsr_reg[3] (.clk (clk), .d (y[21]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[20]));
  CDN_flop \lfsr_reg[4] (.clk (clk), .d (y[22]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[21]));
  CDN_flop \lfsr_reg[5] (.clk (clk), .d (n_3082), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[22]));
  CDN_flop \lfsr_reg[6] (.clk (clk), .d (y[24]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[23]));
  CDN_flop \lfsr_reg[7] (.clk (clk), .d (n_3083), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[24]));
  CDN_flop \lfsr_reg[8] (.clk (clk), .d (y[26]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[25]));
  CDN_flop \lfsr_reg[9] (.clk (clk), .d (y[27]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[26]));
  CDN_flop \lfsr_reg[10] (.clk (clk), .d (n_3084), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[27]));
  CDN_flop \lfsr_reg[11] (.clk (clk), .d (y[17]), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (rst), .srd (1'b0), .q (y[28]));
  CDN_flop round_reg(.clk (clk), .d (1'b0), .sena (1'b0), .aclr (1'b0),
       .apre (1'b0), .srl (n_3118), .srd (n_3086), .q (y[29]));
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
