module task3_top(
    input logic clk,
    input logic rst,

    // Case 1 signals
    output logic rt1,
    output logic rdy1,
    output logic start1,
    output logic endd1,

    // Case 2 signals 
    output logic er2,

    // Case 3 signals 
    output logic er3,
    output logic rdy3,

    // Case 4 signals
    output logic rdy4,
    output logic start4,

    // Case 5 signals
    output logic endd5,
    output logic stop5,
    output logic er5,
    output logic rdy5,
    output logic start5,
    
    // Case 6 signals
    output logic endd6,
    output logic stop6,
    output logic er6,
    output logic rdy6,

    // Case 7 signals
    output logic endd7,
    output logic start7,
    output logic status_valid7,
    output logic instartsv7,

    // Case 8 signals
    output logic rt8,
    output logic enable8,

    // Case 9 signals
    output logic rdy9,
    output logic start9,
    output logic interrupt9,

    // Case 10 singals
    output logic ack10,
    output logic req10
);

    task3_top uufv
    (
        

    );