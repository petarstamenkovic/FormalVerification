bind sv_model black_box_checker c0(.clk(clk), .rst(rst), .x(x), .y(y));

